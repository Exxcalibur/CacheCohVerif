// This RTL design is flattened and obfuscated on purpose.
//start
`include "def.sv"
module  flat_mod_1 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 ,
 parameter TAG_LSB = `TAG_LSB_lv5 , parameter INVALID = 0 )( input rand_rd , input rand_rdx , input randname , input [TAG_MSB : TAG_LSB] tag_randname , input [ASSOC*randname_WID - 1 : 0 ] cache_randname_randname , input [ASSOC*TAG_WID - 1 : 0 ] cache_randname_tag , output reg [ASSOC - 1 : 0 ] access_blk_randname ); integer i; wire [randname_WID - 1 : 0] cache_randname [ASSOC - 1 : 0]; wire [TAG_WID - 1 : 0] cache_tag [ASSOC - 1 : 0]; generate for(genvar gi = 1; gi<=ASSOC; gi++) begin : divide assign cache_randname[gi - 1] = cache_randname_randname[gi*randname_WID - 1 : (gi-1)*randname_WID]; assign cache_tag [gi - 1] = cache_randname_tag [gi*TAG_WID - 1 : (gi-1)*TAG_WID]; end endgenerate always @* begin if(rand_rd || rand_rdx || randname) begin for(i = 0; i < ASSOC; i++) begin if(cache_randname[i] != INVALID && cache_tag[i] == tag_randname) access_blk_randname[i] = 1'b1; else access_blk_randname[i] = 1'b0; end end else begin for(i = 0; i < ASSOC; i++) begin access_blk_randname[i] = 1'b0; end end end endmodule
module  flat_mod_2 #( parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 )( input rand_rd , input rand_rdx , input randname , input [ADDR_WID - 1 : 0] address , output reg [INDEX_MSB : INDEX_LSB] index_randname , output reg [TAG_MSB : TAG_LSB] tag_randname , output reg [OFFSET_MSB : OFFSET_LSB] blk_offset_randname ); reg [ADDR_WID - 1 : 0] zeros = 0; always @ * begin if(rand_rd || rand_rdx || randname) begin index_randname = address[INDEX_MSB : INDEX_LSB]; tag_randname = address[TAG_MSB : TAG_LSB]; blk_offset_randname = address[OFFSET_MSB : OFFSET_LSB]; end else begin index_randname = zeros[INDEX_MSB : INDEX_LSB]; tag_randname = zeros[TAG_MSB : TAG_LSB]; blk_offset_randname = zeros[OFFSET_MSB : OFFSET_LSB]; end end endmodule
module  flat_mod_3 #( parameter ASSOC = `ASSOC_lv5 )( input rand_rd , input rand_rdx , input randname , input [ASSOC - 1 : 0] access_blk_randname , output reg blk_hit_randname ); always @* begin if(rand_rd || rand_rdx || randname) begin if(|access_blk_randname == 1'b1) blk_hit_randname = 1'b1; else blk_hit_randname = 1'b0; end else blk_hit_randname = 1'b0; end endmodule
module blk_to_be_accessed_randname_md #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 )( input blk_hit_randname , input [ASSOC - 1 : 0] access_blk_randname , output reg [ASSOC_WID - 1 : 0] blk_access_randname ); always @* begin blk_access_randname = 0; if(blk_hit_randname) begin for(int i = 0; i < ASSOC; i++) begin if(access_blk_randname[i] == 1'b1) blk_access_randname = i; end end end endmodule
module  flat_mod_4 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 )( input clk , input [1 : 0] core_id , inout [DATA_WID - 1 : 0] data_rand_lv5_lv5 , inout [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 , output lv5_rd , output lv5_wr , input lv5_wr_done , input cpu_rd , input cpu_wr , output cpu_wr_done , inout rand_rd , inout rand_rdx , input rand_lv5_lv5_gnt_randname , output rand_lv5_lv5_req_randname_dl , input rand_lv5_lv5_gnt_randname , output rand_lv5_lv5_req_randname , input [ASSOC_WID - 1 : 0] lru_replacement_randname , output data_in_rand_cpu_lv5_dl , inout data_in_rand_lv5_lv5 , inout randname , input all_invalidation_done , input [randname_WID - 1 : 0] updated_randname_randname , input [randname_WID - 1 : 0] updated_randname_randname , output [randname_WID - 1 : 0] current_randname_randname , output [randname_WID - 1 : 0] current_randname_randname , output shared_local , output cp_in_cache , output invalidation_done , output [ASSOC_WID - 1 : 0] blk_accessed_main ); parameter INVALID = 2'b00; parameter SHARED = 2'b01; parameter EXCLUSIVE = 2'b10; parameter MODIFIED = 2'b11; wire [TAG_MSB : TAG_LSB ] tag_randname; wire [INDEX_MSB : INDEX_LSB ] index_randname; wire [OFFSET_MSB : OFFSET_LSB] blk_offset_randname; wire [TAG_MSB : TAG_LSB ] tag_randname; wire [INDEX_MSB : INDEX_LSB ] index_randname; wire [OFFSET_MSB : OFFSET_LSB] blk_offset_randname; wire [ASSOC*TAG_WID - 1 : 0] cache_randname_tag; wire [ASSOC - 1 : 0] access_blk_randname; wire blk_hit_randname; wire [ASSOC_WID - 1 : 0] blk_access_randname; wire [ASSOC*randname_WID - 1 : 0] cache_randname_randname; wire [ASSOC*randname_WID - 1 : 0] cache_randname_randname; wire [ASSOC*TAG_WID - 1 : 0] cache_randname_tag; wire [ASSOC - 1 : 0] access_blk_randname; wire blk_hit_randname; wire [ASSOC_WID - 1 : 0] blk_access_randname; wire blk_free; wire [ASSOC_WID - 1 : 0] free_blk_num;  flat_mod_20 #( .ASSOC(ASSOC) ) inst_hit_randname_md( .cmd_rd (cpu_rd) , .cmd_wr (cpu_wr) , .access_blk_randname (access_blk_randname) , .blk_hit_randname (blk_hit_randname) );  flat_mod_3 #( .ASSOC(ASSOC) ) inst_hit_randname_md ( .rand_rd (rand_rd), .rand_rdx (rand_rdx), .randname (randname), .access_blk_randname (access_blk_randname), .blk_hit_randname (blk_hit_randname) ); addr_segregator_randname #( .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_addr_segregator_randname ( .cmd_rd (cpu_rd), .cmd_wr (cpu_wr), .address (addr_rand_cpu_lv5), .index_randname (index_randname), .tag_randname (tag_randname), .blk_offset_randname (blk_offset_randname) );  flat_mod_2 #( .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_flat_mod_2 ( .rand_rd (rand_rd), .rand_rdx (rand_rdx), .randname (randname), .address (addr_rand_lv5_lv5), .index_randname (index_randname), .tag_randname (tag_randname), .blk_offset_randname (blk_offset_randname) ); free_blk_md #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .randname_WID(randname_WID), .INVALID(INVALID) ) inst_free_blk_md ( .blk_hit_randname (blk_hit_randname), .cache_randname_randname (cache_randname_randname), .blk_free (blk_free), .free_blk_num (free_blk_num) );  flat_mod_19 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .randname_WID(randname_WID), .TAG_WID(TAG_WID), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .INVALID(INVALID) ) inst_flat_mod_19( .cmd_rd (cpu_rd), .cmd_wr (cpu_wr), .tag_randname (tag_randname), .cache_randname_randname (cache_randname_randname), .cache_randname_tag (cache_randname_tag), .access_blk_randname (access_blk_randname) );  flat_mod_1 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .randname_WID(randname_WID), .TAG_WID(TAG_WID), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .INVALID(INVALID) ) inst_flat_mod_1 ( .rand_rd (rand_rd), .rand_rdx (rand_rdx), .randname (randname), .tag_randname (tag_randname), .cache_randname_randname (cache_randname_randname), .cache_randname_tag (cache_randname_tag), .access_blk_randname (access_blk_randname) ); blk_to_be_accessed_md #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID) ) inst_blk_to_be_accessed_md ( .blk_hit_randname (blk_hit_randname), .access_blk_randname (access_blk_randname), .lru_replacement_randname (lru_replacement_randname), .free_blk_num (free_blk_num), .blk_free (blk_free), .blk_access_randname (blk_access_randname) ); blk_to_be_accessed_randname_md #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID) ) inst_blk_to_be_accessed_randname_md( .blk_hit_randname (blk_hit_randname), .access_blk_randname (access_blk_randname), .blk_access_randname (blk_access_randname) );  flat_mod_11 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .TAG_WID(TAG_WID) ) inst_flat_mod_11 ( .clk (clk), .core_id (core_id), .data_rand_lv5_lv5 (data_rand_lv5_lv5), .addr_rand_lv5_lv5 (addr_rand_lv5_lv5), .data_rand_cpu_lv5 (data_rand_cpu_lv5), .addr_rand_cpu_lv5 (addr_rand_cpu_lv5), .lv5_rd (lv5_rd), .lv5_wr (lv5_wr), .lv5_wr_done (lv5_wr_done), .cpu_rd (cpu_rd), .cpu_wr (cpu_wr), .cpu_wr_done (cpu_wr_done), .rand_rd (rand_rd), .rand_rdx (rand_rdx), .rand_lv5_lv5_gnt_randname (rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname_dl (rand_lv5_lv5_req_randname_dl), .rand_lv5_lv5_gnt_randname (rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname (rand_lv5_lv5_req_randname), .index_randname (index_randname), .index_randname (index_randname), .tag_randname (tag_randname), .tag_randname (tag_randname), .blk_hit_randname (blk_hit_randname), .blk_hit_randname (blk_hit_randname), .blk_free (blk_free), .blk_access_randname (blk_access_randname), .blk_access_randname (blk_access_randname), .lru_replacement_randname (lru_replacement_randname), .data_in_rand_cpu_lv5_dl (data_in_rand_cpu_lv5_dl), .data_in_rand_lv5_lv5 (data_in_rand_lv5_lv5), .randname (randname), .all_invalidation_done (all_invalidation_done), .updated_randname_randname (updated_randname_randname), .updated_randname_randname (updated_randname_randname), .current_randname_randname (current_randname_randname), .current_randname_randname (current_randname_randname), .shared_local (shared_local), .cp_in_cache (cp_in_cache), .invalidation_done (invalidation_done), .blk_accessed_main (blk_accessed_main), .cache_randname_randname (cache_randname_randname), .cache_randname_randname (cache_randname_randname), .cache_randname_tag (cache_randname_tag), .cache_randname_tag (cache_randname_tag) ); endmodule
module  flat_mod_5 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 )( input clk , input [DATA_WID - 1 : 0] data_rand_lv5_lv5 , output [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 , output lv5_rd , input cpu_rd , input rand_lv5_lv5_gnt_randname , output rand_lv5_lv5_req_randname_il , input [ASSOC_WID - 1 : 0] lru_replacement_randname , output data_in_rand_cpu_lv5_il , input data_in_rand_lv5_lv5 , output [ASSOC_WID - 1 : 0] blk_accessed_main ); parameter INVALID = 2'b00; parameter VALID = 2'b01; wire [TAG_MSB : TAG_LSB ] tag_randname; wire [INDEX_MSB : INDEX_LSB ] index_randname; wire [OFFSET_MSB : OFFSET_LSB] blk_offset_randname; wire [ASSOC*randname_WID - 1 : 0] cache_randname_randname; wire [ASSOC*TAG_WID - 1 : 0] cache_randname_tag; wire [ASSOC - 1 : 0] access_blk_randname; wire blk_hit_randname; wire blk_free; wire [ASSOC_WID - 1 : 0] free_blk_num; wire [ASSOC_WID - 1 : 0] blk_access_randname;  flat_mod_20 #( .ASSOC(ASSOC) ) inst_hit_randname_md( .cmd_rd (cpu_rd) , .cmd_wr (1'b0) , .access_blk_randname (access_blk_randname) , .blk_hit_randname (blk_hit_randname) ); addr_segregator_randname #( .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_addr_segregator ( .cmd_rd (cpu_rd), .cmd_wr (1'b0), .address (addr_rand_cpu_lv5), .index_randname (index_randname), .tag_randname (tag_randname), .blk_offset_randname (blk_offset_randname) ); free_blk_md #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .randname_WID(randname_WID), .INVALID(INVALID) ) inst_free_blk_md ( .blk_hit_randname (blk_hit_randname), .cache_randname_randname (cache_randname_randname), .blk_free (blk_free), .free_blk_num (free_blk_num) );  flat_mod_19 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .randname_WID(randname_WID), .TAG_WID(TAG_WID), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .INVALID(INVALID) ) inst_flat_mod_19( .cmd_rd (cpu_rd), .cmd_wr (1'b0), .tag_randname (tag_randname), .cache_randname_randname (cache_randname_randname), .cache_randname_tag (cache_randname_tag), .access_blk_randname (access_blk_randname) ); blk_to_be_accessed_md #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID) ) inst_blk_to_be_accessed_md ( .blk_hit_randname (blk_hit_randname), .access_blk_randname (access_blk_randname), .lru_replacement_randname (lru_replacement_randname), .free_blk_num (free_blk_num), .blk_free (blk_free), .blk_access_randname (blk_access_randname) );  flat_mod_12 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID) ) inst_flat_mod_12( .clk (clk), .data_rand_lv5_lv5 (data_rand_lv5_lv5), .addr_rand_lv5_lv5 (addr_rand_lv5_lv5), .data_rand_cpu_lv5 (data_rand_cpu_lv5), .addr_rand_cpu_lv5 (addr_rand_cpu_lv5), .lv5_rd (lv5_rd), .cpu_rd (cpu_rd), .rand_lv5_lv5_gnt_randname (rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname_il (rand_lv5_lv5_req_randname_il), .index_randname (index_randname), .tag_randname (tag_randname), .blk_hit_randname (blk_hit_randname), .blk_free (blk_free), .blk_access_randname (blk_access_randname), .lru_replacement_randname (lru_replacement_randname), .data_in_rand_cpu_lv5_il (data_in_rand_cpu_lv5_il), .data_in_rand_lv5_lv5 (data_in_rand_lv5_lv5), .blk_accessed_main (blk_accessed_main), .cache_randname_randname (cache_randname_randname), .cache_randname_tag (cache_randname_tag) ); endmodule
module  flat_mod_6 #( parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 )( input [ASSOC_WID - 1 : 0] blk_accessed_main , output [ASSOC_WID - 1 : 0] lru_replacement_randname , input cpu_rd , input cpu_wr , input rand_rd , input rand_rdx , input randname , input shared , input [randname_WID - 1 : 0] current_randname_randname , input [randname_WID - 1 : 0] current_randname_randname , output [randname_WID - 1 : 0] updated_randname_randname , output [randname_WID - 1 : 0] updated_randname_randname , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 ); wire [INDEX_MSB : INDEX_LSB] index_randname; wire [TAG_MSB : TAG_LSB] tag_randname; wire [OFFSET_MSB : OFFSET_LSB] blk_offset_randname;  flat_mod_10 # ( .ASSOC_WID (ASSOC_WID), .INDEX_MSB (INDEX_MSB), .INDEX_LSB (INDEX_LSB), .LRU_VAR_WID (LRU_VAR_WID), .NUM_OF_SETS (NUM_OF_SETS) ) inst_flat_mod_10 ( .index_randname(index_randname), .blk_accessed_main(blk_accessed_main), .lru_replacement_randname(lru_replacement_randname) ); addr_segregator_randname #( .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_addr_segregator ( .cmd_rd (cpu_rd), .cmd_wr (cpu_wr), .address (addr_rand_cpu_lv5), .index_randname (index_randname), .tag_randname (tag_randname), .blk_offset_randname (blk_offset_randname) );  flat_mod_13 #( .randname_WID(randname_WID) ) inst_flat_mod_13 ( .cpu_rd(cpu_rd), .cpu_wr(cpu_wr), .rand_rd(rand_rd), .rand_rdx(rand_rdx), .randname(randname), .shared(shared), .current_randname_randname(current_randname_randname), .current_randname_randname(current_randname_randname), .updated_randname_randname(updated_randname_randname), .updated_randname_randname(updated_randname_randname) ); endmodule
module  flat_mod_7 #( parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 )( input [ASSOC_WID - 1 : 0] blk_accessed_main , output [ASSOC_WID - 1 : 0] lru_replacement_randname , input cpu_rd , input cpu_wr , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 ); wire [INDEX_MSB : INDEX_LSB] index_randname; wire [TAG_MSB : TAG_LSB] tag_randname; wire [OFFSET_MSB : OFFSET_LSB] blk_offset_randname;  flat_mod_10 # ( .ASSOC_WID (ASSOC_WID), .INDEX_MSB (INDEX_MSB), .INDEX_LSB (INDEX_LSB), .LRU_VAR_WID (LRU_VAR_WID), .NUM_OF_SETS (NUM_OF_SETS) ) inst_flat_mod_10 ( .index_randname(index_randname), .blk_accessed_main(blk_accessed_main), .lru_replacement_randname(lru_replacement_randname) ); addr_segregator_randname #( .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_addr_segregator ( .cmd_rd (cpu_rd), .cmd_wr (cpu_wr), .address (addr_rand_cpu_lv5), .index_randname (index_randname), .tag_randname (tag_randname), .blk_offset_randname (blk_offset_randname) ); endmodule
module cache_lv5_multicore #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 , parameter TAG_WID = `TAG_WID_lv5 , parameter IL_DL_ADDR_BOUND = `IL_DL_ADDR_BOUND ) ( input clk , inout [DATA_WID - 1 : 0] data_rand_lv5_lv5 , output [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5_0 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5_0 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5_1 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5_1 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5_2 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5_2 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5_3 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5_3 , output lv5_rd , output lv5_wr , input lv5_wr_done , output cp_in_cache , input [ 3 : 0] cpu_rd , input [ 3 : 0] cpu_wr , output [ 3 : 0] cpu_wr_done , input [ 3 : 0] rand_lv5_lv5_gnt_randname , output [ 3 : 0] rand_lv5_lv5_req_randname , input [ 3 : 0] rand_lv5_lv5_gnt_randname , output [ 3 : 0] rand_lv5_lv5_req_randname , output [ 3 : 0] data_in_rand_cpu_lv5 , inout data_in_rand_lv5_lv5 ); wire [3 : 0] lv5_rd_uni; wire [3 : 0] lv5_wr_uni; wire [3 : 0] cp_in_cache_uni; wire [3 : 0] shared_local; wire shared; wire rand_rd; wire rand_rdx; wire [3 : 0] invalidation_done; wire all_invalidation_done; wire randname; assign lv5_rd = | lv5_rd_uni; assign lv5_wr = | lv5_wr_uni; assign shared = | shared_local; assign all_invalidation_done = | invalidation_done; assign cp_in_cache = | cp_in_cache_uni; cache_lv5_unicore #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .LRU_VAR_WID(LRU_VAR_WID), .NUM_OF_SETS(NUM_OF_SETS), .TAG_WID(TAG_WID), .IL_DL_ADDR_BOUND(IL_DL_ADDR_BOUND) ) inst_cache_lv5_unicore_0 ( .clk(clk), .core_id(0), .data_rand_lv5_lv5(data_rand_lv5_lv5), .addr_rand_lv5_lv5(addr_rand_lv5_lv5), .data_rand_cpu_lv5(data_rand_cpu_lv5_0), .addr_rand_cpu_lv5(addr_rand_cpu_lv5_0), .lv5_rd(lv5_rd_uni[0]), .lv5_wr(lv5_wr_uni[0]), .lv5_wr_done(lv5_wr_done), .cp_in_cache(cp_in_cache_uni[0]), .cpu_rd(cpu_rd[0]), .cpu_wr(cpu_wr[0]), .cpu_wr_done(cpu_wr_done[0]), .rand_rd(rand_rd), .rand_rdx(rand_rdx), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname[0]), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname[0]), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname[0]), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname[0]), .data_in_rand_cpu_lv5(data_in_rand_cpu_lv5[0]), .data_in_rand_lv5_lv5(data_in_rand_lv5_lv5), .randname(randname), .all_invalidation_done(all_invalidation_done), .shared(shared), .shared_local(shared_local[0]), .invalidation_done(invalidation_done[0]) ); cache_lv5_unicore #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .LRU_VAR_WID(LRU_VAR_WID), .NUM_OF_SETS(NUM_OF_SETS), .TAG_WID(TAG_WID), .IL_DL_ADDR_BOUND(IL_DL_ADDR_BOUND) ) inst_cache_lv5_unicore_1 ( .clk(clk), .core_id(1), .data_rand_lv5_lv5(data_rand_lv5_lv5), .addr_rand_lv5_lv5(addr_rand_lv5_lv5), .data_rand_cpu_lv5(data_rand_cpu_lv5_1), .addr_rand_cpu_lv5(addr_rand_cpu_lv5_1), .lv5_rd(lv5_rd_uni[1]), .lv5_wr(lv5_wr_uni[1]), .lv5_wr_done(lv5_wr_done), .cp_in_cache(cp_in_cache_uni[1]), .cpu_rd(cpu_rd[1]), .cpu_wr(cpu_wr[1]), .cpu_wr_done(cpu_wr_done[1]), .rand_rd(rand_rd), .rand_rdx(rand_rdx), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname[1]), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname[1]), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname[1]), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname[1]), .data_in_rand_cpu_lv5(data_in_rand_cpu_lv5[1]), .data_in_rand_lv5_lv5(data_in_rand_lv5_lv5), .randname(randname), .all_invalidation_done(all_invalidation_done), .shared(shared), .shared_local(shared_local[1]), .invalidation_done(invalidation_done[1]) ); cache_lv5_unicore #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .LRU_VAR_WID(LRU_VAR_WID), .NUM_OF_SETS(NUM_OF_SETS), .TAG_WID(TAG_WID), .IL_DL_ADDR_BOUND(IL_DL_ADDR_BOUND) ) inst_cache_lv5_unicore_2 ( .clk(clk), .core_id(2), .data_rand_lv5_lv5(data_rand_lv5_lv5), .addr_rand_lv5_lv5(addr_rand_lv5_lv5), .data_rand_cpu_lv5(data_rand_cpu_lv5_2), .addr_rand_cpu_lv5(addr_rand_cpu_lv5_2), .lv5_rd(lv5_rd_uni[2]), .lv5_wr(lv5_wr_uni[2]), .lv5_wr_done(lv5_wr_done), .cp_in_cache(cp_in_cache_uni[2]), .cpu_rd(cpu_rd[2]), .cpu_wr(cpu_wr[2]), .cpu_wr_done(cpu_wr_done[2]), .rand_rd(rand_rd), .rand_rdx(rand_rdx), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname[2]), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname[2]), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname[2]), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname[2]), .data_in_rand_cpu_lv5(data_in_rand_cpu_lv5[2]), .data_in_rand_lv5_lv5(data_in_rand_lv5_lv5), .randname(randname), .all_invalidation_done(all_invalidation_done), .shared(shared), .shared_local(shared_local[2]), .invalidation_done(invalidation_done[2]) ); cache_lv5_unicore #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .LRU_VAR_WID(LRU_VAR_WID), .NUM_OF_SETS(NUM_OF_SETS), .TAG_WID(TAG_WID), .IL_DL_ADDR_BOUND(IL_DL_ADDR_BOUND) ) inst_cache_lv5_unicore_3 ( .clk(clk), .core_id(3), .data_rand_lv5_lv5(data_rand_lv5_lv5), .addr_rand_lv5_lv5(addr_rand_lv5_lv5), .data_rand_cpu_lv5(data_rand_cpu_lv5_3), .addr_rand_cpu_lv5(addr_rand_cpu_lv5_3), .lv5_rd(lv5_rd_uni[3]), .lv5_wr(lv5_wr_uni[3]), .lv5_wr_done(lv5_wr_done), .cp_in_cache(cp_in_cache_uni[3]), .cpu_rd(cpu_rd[3]), .cpu_wr(cpu_wr[3]), .cpu_wr_done(cpu_wr_done[3]), .rand_rd(rand_rd), .rand_rdx(rand_rdx), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname[3]), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname[3]), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname[3]), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname[3]), .data_in_rand_cpu_lv5(data_in_rand_cpu_lv5[3]), .data_in_rand_lv5_lv5(data_in_rand_lv5_lv5), .randname(randname), .all_invalidation_done(all_invalidation_done), .shared(shared), .shared_local(shared_local[3]), .invalidation_done(invalidation_done[3]) ); endmodule
module cache_lv5_unicore #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 , parameter TAG_WID = `TAG_WID_lv5 , parameter IL_DL_ADDR_BOUND = `IL_DL_ADDR_BOUND )( input clk , input [1 : 0] core_id , inout [DATA_WID - 1 : 0] data_rand_lv5_lv5 , inout [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 , output lv5_rd , output lv5_wr , input lv5_wr_done , input cpu_rd , input cpu_wr , output cpu_wr_done , inout rand_rd , inout rand_rdx , input rand_lv5_lv5_gnt_randname , output rand_lv5_lv5_req_randname , input rand_lv5_lv5_gnt_randname , output rand_lv5_lv5_req_randname , output data_in_rand_cpu_lv5 , inout data_in_rand_lv5_lv5 , inout randname , input all_invalidation_done , input shared , output shared_local , output cp_in_cache , output invalidation_done ); wire cpu_rd_dl; wire cpu_rd_il; wire lv5_rd_dl; wire lv5_rd_il; wire rand_lv5_lv5_req_randname_dl; wire rand_lv5_lv5_req_randname_il; wire data_in_rand_cpu_lv5_dl; wire data_in_rand_cpu_lv5_il; assign cpu_rd_dl = (addr_rand_cpu_lv5 > IL_DL_ADDR_BOUND)? cpu_rd : 1'b0; assign cpu_rd_il = (addr_rand_cpu_lv5 <= IL_DL_ADDR_BOUND)? cpu_rd : 1'b0; assign lv5_rd = lv5_rd_dl | lv5_rd_il; assign rand_lv5_lv5_req_randname = rand_lv5_lv5_req_randname_dl | rand_lv5_lv5_req_randname_il; assign data_in_rand_cpu_lv5 = data_in_rand_cpu_lv5_dl | data_in_rand_cpu_lv5_il;  flat_mod_8 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .LRU_VAR_WID(LRU_VAR_WID), .NUM_OF_SETS(NUM_OF_SETS), .TAG_WID(TAG_WID) ) inst_flat_mod_8 ( .clk(clk), .data_rand_lv5_lv5(data_rand_lv5_lv5), .addr_rand_lv5_lv5(addr_rand_lv5_lv5), .data_rand_cpu_lv5(data_rand_cpu_lv5), .addr_rand_cpu_lv5(addr_rand_cpu_lv5), .lv5_rd(lv5_rd_dl), .lv5_wr(lv5_wr), .lv5_wr_done(lv5_wr_done), .cpu_rd(cpu_rd_dl), .cpu_wr(cpu_wr), .cpu_wr_done(cpu_wr_done), .rand_rd(rand_rd), .rand_rdx(rand_rdx), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname_dl(rand_lv5_lv5_req_randname_dl), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname), .data_in_rand_cpu_lv5_dl(data_in_rand_cpu_lv5_dl), .data_in_rand_lv5_lv5(data_in_rand_lv5_lv5), .randname(randname), .all_invalidation_done(all_invalidation_done), .shared(shared), .shared_local(shared_local), .cp_in_cache(cp_in_cache), .invalidation_done(invalidation_done) );  flat_mod_9 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .LRU_VAR_WID(LRU_VAR_WID), .NUM_OF_SETS(NUM_OF_SETS), .TAG_WID(TAG_WID) ) inst_flat_mod_9 ( .clk(clk), .data_rand_lv5_lv5(data_rand_lv5_lv5), .addr_rand_lv5_lv5(addr_rand_lv5_lv5), .data_rand_cpu_lv5(data_rand_cpu_lv5), .addr_rand_cpu_lv5(addr_rand_cpu_lv5), .lv5_rd(lv5_rd_il), .cpu_rd(cpu_rd_il), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname_il(rand_lv5_lv5_req_randname_il), .data_in_rand_cpu_lv5_il(data_in_rand_cpu_lv5_il), .data_in_rand_lv5_lv5(data_in_rand_lv5_lv5) ); endmodule
module  flat_mod_8 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 , parameter TAG_WID = `TAG_WID_lv5 )( input clk , input [1 : 0] core_id , inout [DATA_WID - 1 : 0] data_rand_lv5_lv5 , inout [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 , output lv5_rd , output lv5_wr , input lv5_wr_done , input cpu_rd , input cpu_wr , output cpu_wr_done , inout rand_rd , inout rand_rdx , input rand_lv5_lv5_gnt_randname , output rand_lv5_lv5_req_randname_dl , input rand_lv5_lv5_gnt_randname , output rand_lv5_lv5_req_randname , output data_in_rand_cpu_lv5_dl , inout data_in_rand_lv5_lv5 , inout randname , input all_invalidation_done , input shared , output shared_local , output cp_in_cache , output invalidation_done ); wire [ASSOC_WID - 1 : 0] lru_replacement_randname; wire [randname_WID - 1 : 0] updated_randname_randname; wire [randname_WID - 1 : 0] updated_randname_randname; wire [ASSOC_WID - 1 : 0] blk_accessed_main; wire [randname_WID - 1 : 0] current_randname_randname; wire [randname_WID - 1 : 0] current_randname_randname;  flat_mod_6 #( .ASSOC_WID(ASSOC_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .LRU_VAR_WID(LRU_VAR_WID), .NUM_OF_SETS(NUM_OF_SETS), .ADDR_WID(ADDR_WID), .randname_WID(randname_WID), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_flat_mod_6 ( .blk_accessed_main(blk_accessed_main), .lru_replacement_randname(lru_replacement_randname), .cpu_rd(cpu_rd), .cpu_wr(cpu_wr), .rand_rd(rand_rd), .rand_rdx(rand_rdx), .randname(randname), .shared(shared), .current_randname_randname(current_randname_randname), .current_randname_randname(current_randname_randname), .updated_randname_randname(updated_randname_randname), .updated_randname_randname(updated_randname_randname), .addr_rand_cpu_lv5(addr_rand_cpu_lv5) );  flat_mod_4 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .TAG_WID(TAG_WID) ) inst_flat_mod_4 ( .clk(clk), .core_id(core_id), .data_rand_lv5_lv5(data_rand_lv5_lv5), .addr_rand_lv5_lv5(addr_rand_lv5_lv5), .data_rand_cpu_lv5(data_rand_cpu_lv5), .addr_rand_cpu_lv5(addr_rand_cpu_lv5), .lv5_rd(lv5_rd), .lv5_wr(lv5_wr), .lv5_wr_done(lv5_wr_done), .cpu_rd(cpu_rd), .cpu_wr(cpu_wr), .cpu_wr_done(cpu_wr_done), .rand_rd(rand_rd), .rand_rdx(rand_rdx), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname_dl(rand_lv5_lv5_req_randname_dl), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname(rand_lv5_lv5_req_randname), .lru_replacement_randname(lru_replacement_randname), .data_in_rand_cpu_lv5_dl(data_in_rand_cpu_lv5_dl), .data_in_rand_lv5_lv5(data_in_rand_lv5_lv5), .randname(randname), .all_invalidation_done(all_invalidation_done), .updated_randname_randname(updated_randname_randname), .updated_randname_randname(updated_randname_randname), .current_randname_randname(current_randname_randname), .current_randname_randname(current_randname_randname), .shared_local(shared_local), .cp_in_cache(cp_in_cache), .invalidation_done(invalidation_done), .blk_accessed_main(blk_accessed_main) );endmodule 
module  flat_mod_9 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 , parameter TAG_WID = `TAG_WID_lv5 )( input clk , input [DATA_WID - 1 : 0] data_rand_lv5_lv5 , output [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 , output lv5_rd , input cpu_rd , input rand_lv5_lv5_gnt_randname , output rand_lv5_lv5_req_randname_il , output data_in_rand_cpu_lv5_il , input data_in_rand_lv5_lv5 ); wire [ASSOC_WID - 1 : 0] lru_replacement_randname; wire [ASSOC_WID - 1 : 0] blk_accessed_main;  flat_mod_7 #( .ASSOC_WID(ASSOC_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .LRU_VAR_WID(LRU_VAR_WID), .NUM_OF_SETS(NUM_OF_SETS), .ADDR_WID(ADDR_WID), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_flat_mod_7 ( .blk_accessed_main(blk_accessed_main), .lru_replacement_randname(lru_replacement_randname), .cpu_rd(cpu_rd), .cpu_wr(1'b0), .addr_rand_cpu_lv5(addr_rand_cpu_lv5) );  flat_mod_5 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID), .TAG_WID(TAG_WID) ) inst_flat_mod_5 ( .clk(clk), .data_rand_lv5_lv5(data_rand_lv5_lv5), .addr_rand_lv5_lv5(addr_rand_lv5_lv5), .data_rand_cpu_lv5(data_rand_cpu_lv5), .addr_rand_cpu_lv5(addr_rand_cpu_lv5), .lv5_rd(lv5_rd), .cpu_rd(cpu_rd), .rand_lv5_lv5_gnt_randname(rand_lv5_lv5_gnt_randname), .rand_lv5_lv5_req_randname_il(rand_lv5_lv5_req_randname_il), .lru_replacement_randname(lru_replacement_randname), .data_in_rand_cpu_lv5_il(data_in_rand_cpu_lv5_il), .data_in_rand_lv5_lv5(data_in_rand_lv5_lv5), .blk_accessed_main(blk_accessed_main) ); endmodule
module  flat_mod_10 #( parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 ) ( input [INDEX_MSB : INDEX_LSB ] index_randname , input [ASSOC_WID - 1 : 0 ] blk_accessed_main , output reg [ASSOC_WID - 1 : 0 ] lru_replacement_randname ); parameter BLK0_REPLACEMENT = 3'b00x; parameter BLK1_REPLACEMENT = 3'b01x; parameter BLK2_REPLACEMENT = 3'b1x0; parameter BLK3_REPLACEMENT = 3'b1x1; reg [LRU_VAR_WID - 1 : 0] lru_var [NUM_OF_SETS - 1 : 0]; always @ * begin casex (lru_var[index_randname]) BLK0_REPLACEMENT: lru_replacement_randname = 2'b00; BLK1_REPLACEMENT: lru_replacement_randname = 2'b01; BLK2_REPLACEMENT: lru_replacement_randname = 2'b10; BLK3_REPLACEMENT: lru_replacement_randname = 2'b11; default: lru_replacement_randname = 2'b00; endcase end always @ * begin case (blk_accessed_main) 3'b000: begin lru_var[index_randname][2:1] = 2'b11; end 3'b001: begin lru_var[index_randname][2:1] = 2'b10; end 3'b010: begin lru_var[index_randname][2] = 1'b0; lru_var[index_randname][0] = 1'b1; end 3'b011: begin lru_var[index_randname][2] = 1'b0; lru_var[index_randname][0] = 1'b0; end default: lru_var[index_randname] = 3'b0; endcase end endmodule
module  flat_mod_11 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 )( input clk , input [1 : 0] core_id , inout [DATA_WID - 1 : 0] data_rand_lv5_lv5 , inout [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 , output reg lv5_rd , output reg lv5_wr , input lv5_wr_done , input cpu_rd , input cpu_wr , output reg cpu_wr_done , inout rand_rd , inout rand_rdx , input rand_lv5_lv5_gnt_randname , output reg rand_lv5_lv5_req_randname_dl , input rand_lv5_lv5_gnt_randname , output reg rand_lv5_lv5_req_randname , input [INDEX_MSB : INDEX_LSB] index_randname , input [INDEX_MSB : INDEX_LSB] index_randname , input [TAG_MSB : TAG_LSB] tag_randname , input [TAG_MSB : TAG_LSB] tag_randname , input blk_hit_randname , input blk_hit_randname , input blk_free , input [ASSOC_WID - 1 : 0] blk_access_randname , input [ASSOC_WID - 1 : 0] blk_access_randname , input [ASSOC_WID - 1 : 0] lru_replacement_randname , output reg data_in_rand_cpu_lv5_dl , inout data_in_rand_lv5_lv5 , inout randname , input all_invalidation_done , input [randname_WID - 1 : 0] updated_randname_randname , input [randname_WID - 1 : 0] updated_randname_randname , output [randname_WID - 1 : 0] current_randname_randname , output [randname_WID - 1 : 0] current_randname_randname , output reg shared_local , output reg cp_in_cache , output reg invalidation_done , output reg [ASSOC_WID - 1 : 0] blk_accessed_main , output reg [ASSOC*randname_WID - 1 : 0] cache_randname_randname , output reg [ASSOC*randname_WID - 1 : 0] cache_randname_randname , output reg [ASSOC*TAG_WID - 1 : 0] cache_randname_tag , output reg [ASSOC*TAG_WID - 1 : 0] cache_randname_tag ); parameter INVALID = 2'b00; parameter SHARED = 2'b01; parameter EXCLUSIVE = 2'b10; parameter MODIFIED = 2'b11; reg [CACHE_DATA_WID - 1 : 0] cache_var [0 : CACHE_DEPTH - 1]; reg [CACHE_TAG_randname_WID - 1 : 0] cache_randname_contr [0 : CACHE_DEPTH - 1]; reg [DATA_WID - 1 : 0] data_rand_lv5_lv5_reg; reg [ADDR_WID - 1 : 0] addr_rand_lv5_lv5_reg; reg [DATA_WID - 1 : 0] data_rand_cpu_lv5_reg; reg data_in_rand_lv5_lv5_reg; reg rand_rd_reg; reg rand_rdx_reg; reg randname_reg; initial begin for (int i = 0; i<CACHE_DEPTH; i++) begin cache_var[i] = {CACHE_DATA_WID{1'b0}}; cache_randname_contr[i] = {CACHE_TAG_randname_WID{1'b0}}; end end assign data_rand_lv5_lv5 = data_rand_lv5_lv5_reg; assign addr_rand_lv5_lv5 = addr_rand_lv5_lv5_reg; assign data_rand_cpu_lv5 = data_rand_cpu_lv5_reg; assign data_in_rand_lv5_lv5 = data_in_rand_lv5_lv5_reg; assign rand_rd = rand_rd_reg; assign rand_rdx = rand_rdx_reg; assign randname = randname_reg; generate for(genvar gi = 1; gi<=ASSOC; gi++) begin assign cache_randname_randname [gi*randname_WID - 1 : (gi-1)*randname_WID] = cache_randname_contr[{index_randname,{ASSOC_WID{1'b0}}}+gi-1][CACHE_randname_MSB : CACHE_randname_LSB]; assign cache_randname_tag [gi*TAG_WID - 1 : (gi-1)*TAG_WID ] = cache_randname_contr[{index_randname,{ASSOC_WID{1'b0}}}+gi-1][CACHE_TAG_MSB : CACHE_TAG_LSB ]; assign cache_randname_randname[gi*randname_WID - 1 : (gi-1)*randname_WID] = cache_randname_contr[{index_randname,{ASSOC_WID{1'b0}}}+gi-1][CACHE_randname_MSB : CACHE_randname_LSB]; assign cache_randname_tag [gi*TAG_WID - 1 : (gi-1)*TAG_WID ] = cache_randname_contr[{index_randname,{ASSOC_WID{1'b0}}}+gi-1][CACHE_TAG_MSB : CACHE_TAG_LSB ]; end endgenerate assign current_randname_randname = `CACHE_CURRENT_randname_randname; assign current_randname_randname = `CACHE_CURRENT_randname_randname; always @(posedge clk) begin data_rand_cpu_lv5_reg <= 32'hz; data_rand_lv5_lv5_reg <= 32'hz; addr_rand_lv5_lv5_reg <= 32'hz; rand_rd_reg <= 1'bz; rand_rdx_reg <= 1'bz; data_in_rand_lv5_lv5_reg <= 1'bz; randname_reg <= 1'bz; invalidation_done <= 1'b0; rand_lv5_lv5_req_randname_dl <= 1'b0; rand_lv5_lv5_req_randname <= 1'b0; data_in_rand_cpu_lv5_dl <= 1'b0; lv5_rd <= 1'b0; lv5_wr <= 1'b0; shared_local <= 1'b0; cpu_wr_done <= 1'b0; cp_in_cache <= 1'b0; if(cpu_rd && blk_hit_randname) begin data_rand_cpu_lv5_reg <= cache_var[{index_randname,blk_access_randname}]; data_in_rand_cpu_lv5_dl <= 1'b1; blk_accessed_main <= blk_access_randname; end else if(cpu_rd && !blk_hit_randname) begin rand_lv5_lv5_req_randname_dl <= 1'b1; if(blk_free) begin if(rand_lv5_lv5_gnt_randname) begin rand_rd_reg <= 1'b1; lv5_rd <= 1'b1; addr_rand_lv5_lv5_reg <= {tag_randname, index_randname, 2'b00}; if(data_in_rand_lv5_lv5) begin if(updated_randname_randname == SHARED) cache_var[{index_randname,blk_access_randname}] <= data_rand_lv5_lv5; else cache_var[{index_randname,blk_access_randname}] <= {tag_randname, index_randname, 2'b00}; `CACHE_CURRENT_randname_randname <= updated_randname_randname; `CACHE_CURRENT_TAG_randname <= tag_randname; rand_lv5_lv5_req_randname_dl <= 1'b0; rand_rd_reg <= 1'bz; lv5_rd <= 1'b0; addr_rand_lv5_lv5_reg <= 32'hz; end end end else if(!blk_free) begin case (`CACHE_CURRENT_randname_randname) SHARED: `CACHE_CURRENT_randname_randname <= INVALID; EXCLUSIVE: `CACHE_CURRENT_randname_randname <= INVALID; MODIFIED: begin if(rand_lv5_lv5_gnt_randname) begin addr_rand_lv5_lv5_reg <= {`CACHE_CURRENT_TAG_randname,index_randname,2'b00}; lv5_wr <= 1'b1; data_rand_lv5_lv5_reg <= cache_var[{index_randname,blk_access_randname}]; if(lv5_wr_done) begin `CACHE_CURRENT_randname_randname <= INVALID; addr_rand_lv5_lv5_reg <= 32'hz; lv5_wr <= 1'b0; data_rand_lv5_lv5_reg <= 32'hz; end end end default: `CACHE_CURRENT_randname_randname <= INVALID; endcase end end if(cpu_wr) begin rand_lv5_lv5_req_randname_dl <= 1'b1; if(blk_hit_randname) begin case (`CACHE_CURRENT_randname_randname) SHARED: begin if(rand_lv5_lv5_gnt_randname) begin randname_reg <= 1'b1; addr_rand_lv5_lv5_reg <= {tag_randname,index_randname,2'b00}; if(all_invalidation_done) begin cache_var[{index_randname,blk_access_randname}] <= data_rand_cpu_lv5; `CACHE_CURRENT_randname_randname <= updated_randname_randname; cpu_wr_done <= 1'b1; blk_accessed_main <= blk_access_randname; rand_lv5_lv5_req_randname_dl <= 1'b0; randname_reg <= 1'bz; addr_rand_lv5_lv5_reg <= 32'hz; end end end default: begin cache_var[{index_randname,blk_access_randname}] <= data_rand_cpu_lv5; `CACHE_CURRENT_randname_randname <= updated_randname_randname; cpu_wr_done <= 1'b1; blk_accessed_main <= blk_access_randname; rand_lv5_lv5_req_randname_dl <= 1'b0; end endcase end else if (blk_free) begin if(rand_lv5_lv5_gnt_randname) begin rand_rdx_reg <= 1'b1; lv5_rd <= 1'b1; addr_rand_lv5_lv5_reg <= {tag_randname,index_randname,2'b00}; if(data_in_rand_lv5_lv5) begin cache_var[{index_randname,blk_access_randname}] <= data_rand_lv5_lv5; `CACHE_CURRENT_randname_randname <= updated_randname_randname; `CACHE_CURRENT_TAG_randname <= tag_randname; rand_lv5_lv5_req_randname_dl <= 1'b0; rand_rdx_reg <= 1'b0; lv5_rd <= 1'b0; addr_rand_lv5_lv5_reg <= 32'hz; end end end else begin case (`CACHE_CURRENT_randname_randname) SHARED: `CACHE_CURRENT_randname_randname <= INVALID; EXCLUSIVE: `CACHE_CURRENT_randname_randname <= INVALID; MODIFIED: begin if(rand_lv5_lv5_gnt_randname) begin addr_rand_lv5_lv5_reg <= {`CACHE_CURRENT_TAG_randname,index_randname,2'b00}; lv5_wr <= 1'b1; data_rand_lv5_lv5_reg <= cache_var[{index_randname,blk_access_randname}]; if(lv5_wr_done) begin `CACHE_CURRENT_randname_randname <= INVALID; addr_rand_lv5_lv5_reg <= 32'hz; lv5_wr <= 1'b0; data_rand_lv5_lv5_reg <= 32'hz; end end end default: `CACHE_CURRENT_randname_randname <= INVALID; endcase end end if(blk_hit_randname && (rand_lv5_lv5_gnt_randname != 1'b1)) begin if(randname) begin shared_local <= 1'b1; invalidation_done <= 1'b1; end else if(rand_rdx) begin cp_in_cache <= 1'b1; case (`CACHE_CURRENT_randname_randname) SHARED: begin shared_local <= 1'b1; `CACHE_CURRENT_randname_randname <= updated_randname_randname; end MODIFIED: begin rand_lv5_lv5_req_randname <= 1'b1; if(rand_lv5_lv5_gnt_randname) begin data_rand_lv5_lv5_reg <= cache_var[{index_randname,blk_access_randname}]; lv5_wr <= 1'b1; if(lv5_wr_done) begin `CACHE_CURRENT_randname_randname <= updated_randname_randname; lv5_wr <= 1'b0; data_rand_lv5_lv5_reg <= 32'hz; end end end default: `CACHE_CURRENT_randname_randname <= updated_randname_randname; endcase end else if(rand_rd) begin rand_lv5_lv5_req_randname <= 1'b1; cp_in_cache <= 1'b1; if(data_in_rand_lv5_lv5 && !rand_lv5_lv5_gnt_randname) rand_lv5_lv5_req_randname <= 1'b0; if(rand_lv5_lv5_gnt_randname) begin case (`CACHE_CURRENT_randname_randname) MODIFIED: begin data_rand_lv5_lv5_reg <= cache_var[{index_randname,blk_access_randname}]; lv5_wr <= 1'b1; if(lv5_wr_done) begin data_in_rand_lv5_lv5_reg <= 1'b1; shared_local <= 1'b1; `CACHE_CURRENT_randname_randname <= updated_randname_randname; lv5_wr <= 1'b0; end end default: begin data_rand_lv5_lv5_reg <= cache_var[{index_randname,blk_access_randname}]; data_in_rand_lv5_lv5_reg <= 1'b1; shared_local <= 1'b1; `CACHE_CURRENT_randname_randname <= updated_randname_randname; end endcase end end end end endmodule
module  flat_mod_12 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 )( input clk , input [DATA_WID - 1 : 0] data_rand_lv5_lv5 , output reg [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_cpu_lv5 , input [ADDR_WID - 1 : 0] addr_rand_cpu_lv5 , output reg lv5_rd , input cpu_rd , input rand_lv5_lv5_gnt_randname , output reg rand_lv5_lv5_req_randname_il , input [INDEX_MSB : INDEX_LSB] index_randname , input [TAG_MSB : TAG_LSB] tag_randname , input blk_hit_randname , input blk_free , input [ASSOC_WID - 1 : 0] blk_access_randname , input [ASSOC_WID - 1 : 0] lru_replacement_randname , output reg data_in_rand_cpu_lv5_il , input data_in_rand_lv5_lv5 , output reg [ASSOC_WID - 1 : 0] blk_accessed_main , output reg [ASSOC*randname_WID - 1 : 0] cache_randname_randname , output reg [ASSOC*TAG_WID - 1 : 0] cache_randname_tag ); integer i; parameter INVALID = 2'b00; parameter VALID = 2'b01; reg [CACHE_DATA_WID - 1 : 0] cache_var [0 : CACHE_DEPTH - 1]; reg [CACHE_TAG_randname_WID - 1 : 0] cache_randname_contr [0 : CACHE_DEPTH - 1]; reg [DATA_WID - 1 : 0] data_rand_cpu_lv5_reg; reg [31:0] zeros = 32'h0; initial begin for (i = 0; i<CACHE_DEPTH; i++) begin cache_var[i] = {CACHE_DATA_WID{1'b0}}; cache_randname_contr[i] = {CACHE_TAG_randname_WID{1'b0}}; end end assign data_rand_cpu_lv5 = data_rand_cpu_lv5_reg; generate for(genvar gi = 1; gi<=ASSOC; gi++) begin assign cache_randname_randname[gi*randname_WID - 1 : (gi-1)*randname_WID] = cache_randname_contr[{index_randname,{ASSOC_WID{1'b0}}}+gi-1][CACHE_randname_MSB : CACHE_randname_LSB]; assign cache_randname_tag [gi*TAG_WID - 1 : (gi-1)*TAG_WID ] = cache_randname_contr[{index_randname,{ASSOC_WID{1'b0}}}+gi-1][CACHE_TAG_MSB : CACHE_TAG_LSB ]; end endgenerate always @(posedge clk) begin data_rand_cpu_lv5_reg <= 32'hz; rand_lv5_lv5_req_randname_il <= 1'b0; data_in_rand_cpu_lv5_il <= 1'b0; lv5_rd <= 1'b0; addr_rand_lv5_lv5 <= 32'hz; if(cpu_rd) begin if(blk_hit_randname) begin data_rand_cpu_lv5_reg <= cache_var[{index_randname,blk_access_randname}]; data_in_rand_cpu_lv5_il <= 1'b1; blk_accessed_main <= blk_access_randname; end else if(blk_free) begin rand_lv5_lv5_req_randname_il <= 1'b1; if(rand_lv5_lv5_gnt_randname) begin lv5_rd <= 1'b1; addr_rand_lv5_lv5 <= {tag_randname, index_randname, {OFFSET_WID{1'b0}}}; if(data_in_rand_lv5_lv5) begin cache_var[{index_randname,blk_access_randname}] <= data_rand_lv5_lv5; `CACHE_CURRENT_randname <= VALID; `CACHE_CURRENT_TAG <= tag_randname; rand_lv5_lv5_req_randname_il <= 1'b0; lv5_rd <= 1'b0; addr_rand_lv5_lv5 <= 32'hz; end end end else begin `CACHE_CURRENT_randname <= INVALID; end end end endmodule
module  flat_mod_13 #( parameter randname_WID = `randname_WID_lv5 )( input cpu_rd , input cpu_wr , input rand_rd , input rand_rdx , input randname , input shared , input [randname_WID - 1 : 0] current_randname_randname , input [randname_WID - 1 : 0] current_randname_randname , output reg [randname_WID - 1 : 0] updated_randname_randname , output reg [randname_WID - 1 : 0] updated_randname_randname ); parameter INVALID = 2'b00; parameter SHARED = 2'b01; parameter EXCLUSIVE = 2'b10; parameter MODIFIED = 2'b11; always @* begin updated_randname_randname = INVALID; case (current_randname_randname) MODIFIED: begin updated_randname_randname = MODIFIED; end EXCLUSIVE: begin if (cpu_rd) updated_randname_randname = EXCLUSIVE; else if (cpu_wr) updated_randname_randname = MODIFIED; else updated_randname_randname = EXCLUSIVE; end SHARED: begin if (cpu_rd) updated_randname_randname = SHARED; else if (cpu_wr) updated_randname_randname = MODIFIED; else updated_randname_randname = SHARED; end INVALID: begin if (cpu_rd && !shared) updated_randname_randname = EXCLUSIVE; else if (cpu_rd && shared) updated_randname_randname = SHARED; else if (cpu_wr) updated_randname_randname = MODIFIED; else updated_randname_randname = INVALID; end default: updated_randname_randname = INVALID; endcase end always @* begin updated_randname_randname = INVALID; case(current_randname_randname) MODIFIED: begin if(rand_rd) updated_randname_randname = SHARED; else if(rand_rdx) updated_randname_randname = INVALID; else updated_randname_randname = MODIFIED; end EXCLUSIVE: begin if(rand_rd) updated_randname_randname = SHARED; else if(rand_rdx) updated_randname_randname = INVALID; else updated_randname_randname = EXCLUSIVE; end SHARED: begin if(rand_rdx || randname) updated_randname_randname = INVALID; else updated_randname_randname = SHARED; end INVALID: begin updated_randname_randname = INVALID; end default: updated_randname_randname = INVALID; endcase end endmodule
module  flat_mod_14 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 )( input clk , input [ASSOC_WID - 1 : 0] lru_replacement_randname , output [ASSOC_WID - 1 : 0] blk_accessed_main , inout [DATA_WID - 1 : 0] data_rand_lv5_lv5 , input [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_lv5_mem , output [ADDR_WID - 1 : 0] addr_rand_lv5_mem , output mem_rd , output mem_wr , input mem_wr_done , input lv5_rd , input lv5_wr , output lv5_wr_done , input cp_in_cache , input rand_lv5_lv5_gnt_lv5 , output rand_lv5_lv5_req_lv5 , output data_in_rand_lv5_lv5 , input data_in_rand_lv5_mem ); parameter INVALID = 2'b00; parameter VALID = 2'b01; parameter MODIFIED = 2'b10; wire [TAG_MSB : TAG_LSB ] tag_randname;
  wire [INDEX_MSB : INDEX_LSB ] index_randname; wire [OFFSET_MSB : OFFSET_LSB] blk_offset_randname; wire [ASSOC*randname_WID - 1 : 0] cache_randname_randname; wire [ASSOC*TAG_WID - 1 : 0] cache_randname_tag; wire [ASSOC - 1 : 0] access_blk_randname; wire blk_hit_randname; wire blk_free; wire [ASSOC_WID - 1 : 0] free_blk_num; wire [ASSOC_WID - 1 : 0] blk_access_randname; 
  flat_mod_20 #( .ASSOC(ASSOC) ) inst_hit_randname_md( .cmd_rd (lv5_rd) , .cmd_wr (lv5_wr) , .access_blk_randname (access_blk_randname) , .blk_hit_randname (blk_hit_randname) ); addr_segregator_randname #( .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_addr_segregator ( .cmd_rd (lv5_rd), .cmd_wr (lv5_wr), .address (addr_rand_lv5_lv5), .index_randname (index_randname), .tag_randname (tag_randname), .blk_offset_randname (blk_offset_randname) ); free_blk_md #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .randname_WID(randname_WID), .INVALID(INVALID) ) inst_free_blk_md ( .blk_hit_randname (blk_hit_randname), .cache_randname_randname (cache_randname_randname), .blk_free (blk_free), .free_blk_num (free_blk_num) ); 
   flat_mod_19 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .randname_WID(randname_WID), .TAG_WID(TAG_WID), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .INVALID(INVALID) ) inst_blk_randname_md( .cmd_rd (lv5_rd), .cmd_wr (lv5_wr), .tag_randname (tag_randname), .cache_randname_randname (cache_randname_randname), .cache_randname_tag (cache_randname_tag), .access_blk_randname (access_blk_randname) ); 
  blk_to_be_accessed_md #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID) ) inst_blk_to_be_accessed_md ( .blk_hit_randname (blk_hit_randname), .access_blk_randname (access_blk_randname), .lru_replacement_randname (lru_replacement_randname), .free_blk_num (free_blk_num), .blk_free (blk_free), .blk_access_randname (blk_access_randname) );
   flat_mod_18 #( .ASSOC(ASSOC), .ASSOC_WID(ASSOC_WID), .DATA_WID(DATA_WID), .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB), .CACHE_DATA_WID(CACHE_DATA_WID), .CACHE_TAG_MSB(CACHE_TAG_MSB), .CACHE_TAG_LSB(CACHE_TAG_LSB), .CACHE_DEPTH(CACHE_DEPTH), .CACHE_randname_MSB(CACHE_randname_MSB), .CACHE_randname_LSB(CACHE_randname_LSB), .CACHE_TAG_randname_WID(CACHE_TAG_randname_WID), .randname_WID(randname_WID), .OFFSET_WID(OFFSET_WID) ) inst_flat_mod_18( .clk (clk), .data_rand_lv5_lv5 (data_rand_lv5_lv5), .addr_rand_lv5_lv5 (addr_rand_lv5_lv5), .data_rand_lv5_mem (data_rand_lv5_mem), .addr_rand_lv5_mem (addr_rand_lv5_mem), .mem_rd (mem_rd), .mem_wr (mem_wr), .mem_wr_done (mem_wr_done), .lv5_rd (lv5_rd), .lv5_wr (lv5_wr), .lv5_wr_done (lv5_wr_done), .cp_in_cache (cp_in_cache), .rand_lv5_lv5_gnt_lv5 (rand_lv5_lv5_gnt_lv5), .rand_lv5_lv5_req_lv5 (rand_lv5_lv5_req_lv5), .index_randname (index_randname), .tag_randname (tag_randname), .blk_hit_randname (blk_hit_randname), .blk_free (blk_free), .blk_access_randname (blk_access_randname), .lru_replacement_randname (lru_replacement_randname), .data_in_rand_lv5_lv5 (data_in_rand_lv5_lv5), .data_in_rand_lv5_mem (data_in_rand_lv5_mem), .blk_accessed_main (blk_accessed_main), .cache_randname_randname (cache_randname_randname), .cache_randname_tag (cache_randname_tag) ); endmodule
module  flat_mod_15 #( parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 )( input [ASSOC_WID - 1 : 0] blk_accessed_main , output [ASSOC_WID - 1 : 0] lru_replacement_randname , input lv5_rd , input lv5_wr , input [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 ); wire [INDEX_MSB : INDEX_LSB] index_randname;
wire [TAG_MSB : TAG_LSB] tag_randname; wire [OFFSET_MSB : OFFSET_LSB] blk_offset_randname;  flat_mod_17 # ( .ASSOC_WID (ASSOC_WID), .INDEX_MSB (INDEX_MSB), .INDEX_LSB (INDEX_LSB), .LRU_VAR_WID (LRU_VAR_WID), .NUM_OF_SETS (NUM_OF_SETS) ) inst_flat_mod_17 ( .index_randname(index_randname), .blk_accessed_main(blk_accessed_main), .lru_replacement_randname(lru_replacement_randname) ); addr_segregator_randname #( .ADDR_WID(ADDR_WID), .INDEX_MSB(INDEX_MSB), .INDEX_LSB(INDEX_LSB), .OFFSET_MSB(OFFSET_MSB), .OFFSET_LSB(OFFSET_LSB), .TAG_MSB(TAG_MSB), .TAG_LSB(TAG_LSB) ) inst_addr_segregator ( .cmd_rd (lv5_rd), .cmd_wr (lv5_wr), .address (addr_rand_lv5_lv5), .index_randname (index_randname), .tag_randname (tag_randname), .blk_offset_randname (blk_offset_randname) ); endmodule
 module  flat_mod_16 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 ) ( input clk , inout [DATA_WID - 1 : 0] data_rand_lv5_lv5 , input [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_lv5_mem , output [ADDR_WID - 1 : 0] addr_rand_lv5_mem , output mem_rd , output mem_wr , input mem_wr_done , input lv5_rd , input lv5_wr , output lv5_wr_done , input cp_in_cache , input rand_lv5_lv5_gnt_lv5 , output rand_lv5_lv5_req_lv5 , output data_in_rand_lv5_lv5 , input data_in_rand_lv5_mem ); wire [ASSOC_WID - 1 : 0] lru_replacement_randname ; wire [ASSOC_WID - 1 : 0] blk_accessed_main ;  flat_mod_14 inst_flat_mod_14 ( .clk (clk), .lru_replacement_randname (lru_replacement_randname), .blk_accessed_main (blk_accessed_main), .data_rand_lv5_lv5 (data_rand_lv5_lv5), .addr_rand_lv5_lv5 (addr_rand_lv5_lv5), .data_rand_lv5_mem (data_rand_lv5_mem), .addr_rand_lv5_mem (addr_rand_lv5_mem), .mem_rd (mem_rd), .mem_wr (mem_wr), .mem_wr_done (mem_wr_done), .lv5_rd (lv5_rd), .lv5_wr (lv5_wr), .lv5_wr_done (lv5_wr_done), .cp_in_cache (cp_in_cache), .rand_lv5_lv5_gnt_lv5 (rand_lv5_lv5_gnt_lv5), .rand_lv5_lv5_req_lv5 (rand_lv5_lv5_req_lv5), .data_in_rand_lv5_lv5 (data_in_rand_lv5_lv5), .data_in_rand_lv5_mem (data_in_rand_lv5_mem) );  flat_mod_15 inst_flat_mod_15 ( .blk_accessed_main (blk_accessed_main), .lru_replacement_randname (lru_replacement_randname), .lv5_rd (lv5_rd), .lv5_wr (lv5_wr), .addr_rand_lv5_lv5 (addr_rand_lv5_lv5) );endmodule
module  flat_mod_17 #( parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter LRU_VAR_WID = `LRU_VAR_WID_lv5 , parameter NUM_OF_SETS = `NUM_OF_SETS_lv5 ) ( input [INDEX_MSB : INDEX_LSB ] index_randname , input [ASSOC_WID - 1 : 0 ] blk_accessed_main , output reg [ASSOC_WID - 1 : 0 ] lru_replacement_randname ); parameter BLK0_REPLACEMENT = 7'b00x0xxx; parameter BLK1_REPLACEMENT = 7'b00x1xxx; parameter BLK2_REPLACEMENT = 7'b01xx0xx; parameter BLK3_REPLACEMENT = 7'b01xx1xx; parameter BLK4_REPLACEMENT = 7'b1x0xx0x; parameter BLK5_REPLACEMENT = 7'b1x0xx1x; parameter BLK6_REPLACEMENT = 7'b1x1xxx0; parameter BLK7_REPLACEMENT = 7'b1x1xxx1; reg [LRU_VAR_WID - 1 : 0] lru_var [NUM_OF_SETS - 1 : 0]; always @ * begin casex (lru_var[index_randname]) BLK0_REPLACEMENT: lru_replacement_randname = 3'b000; BLK1_REPLACEMENT: lru_replacement_randname = 3'b001; BLK2_REPLACEMENT: lru_replacement_randname = 3'b010; BLK3_REPLACEMENT: lru_replacement_randname = 3'b011; BLK4_REPLACEMENT: lru_replacement_randname = 3'b100; BLK5_REPLACEMENT: lru_replacement_randname = 3'b101; BLK6_REPLACEMENT: lru_replacement_randname = 3'b110; BLK7_REPLACEMENT: lru_replacement_randname = 3'b111; default: lru_replacement_randname = 3'b000; endcase end always @ * begin case (blk_accessed_main) 3'b000: begin lru_var[index_randname][6:5] = 2'b11; lru_var[index_randname][3] = 1'b1; end 3'b001: begin lru_var[index_randname][6:5] = 2'b11; lru_var[index_randname][3] = 1'b0; end 3'b010: begin lru_var[index_randname][6:5] = 2'b10; lru_var[index_randname][2] = 1'b1; end 3'b011: begin lru_var[index_randname][6:5] = 2'b10; lru_var[index_randname][2] = 1'b0; end 3'b100: begin lru_var[index_randname][6] = 1'b0; lru_var[index_randname][4] = 1'b1; lru_var[index_randname][1] = 1'b1; end 3'b101: begin lru_var[index_randname][6] = 1'b0; lru_var[index_randname][4] = 1'b1; lru_var[index_randname][1] = 1'b0; end 3'b110: begin lru_var[index_randname][6] = 1'b0; lru_var[index_randname][4] = 1'b0; lru_var[index_randname][0] = 1'b1; end 3'b111: begin lru_var[index_randname][6] = 1'b0; lru_var[index_randname][4] = 1'b0; lru_var[index_randname][0] = 1'b0; end default: lru_var[index_randname] = 7'b0; endcase end endmodule 
module  flat_mod_18 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter DATA_WID = `DATA_WID_lv5 , parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter CACHE_DATA_WID = `CACHE_DATA_WID_lv5 , parameter CACHE_TAG_MSB = `CACHE_TAG_MSB_lv5 , parameter CACHE_TAG_LSB = `CACHE_TAG_LSB_lv5 , parameter CACHE_DEPTH = `CACHE_DEPTH_lv5 , parameter CACHE_randname_MSB = `CACHE_randname_MSB_lv5 , parameter CACHE_randname_LSB = `CACHE_randname_LSB_lv5 , parameter CACHE_TAG_randname_WID = `CACHE_TAG_randname_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter OFFSET_WID = `OFFSET_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 )( input clk , inout [DATA_WID - 1 : 0] data_rand_lv5_lv5 , input [ADDR_WID - 1 : 0] addr_rand_lv5_lv5 , inout [DATA_WID - 1 : 0] data_rand_lv5_mem , output reg [ADDR_WID - 1 : 0] addr_rand_lv5_mem , output reg mem_rd , output reg mem_wr , input mem_wr_done , input lv5_rd , input lv5_wr , output reg lv5_wr_done , input cp_in_cache , input rand_lv5_lv5_gnt_lv5 , output reg rand_lv5_lv5_req_lv5 ,
input [INDEX_MSB : INDEX_LSB] index_randname , input [TAG_MSB : TAG_LSB] tag_randname , input blk_hit_randname , input blk_free , input [ASSOC_WID - 1 : 0] blk_access_randname , input [ASSOC_WID - 1 : 0] lru_replacement_randname , output reg data_in_rand_lv5_lv5 , input data_in_rand_lv5_mem , output reg [ASSOC_WID - 1 : 0] blk_accessed_main , output reg [ASSOC*randname_WID - 1 : 0] cache_randname_randname , output reg [ASSOC*TAG_WID - 1 : 0] cache_randname_tag ); integer i; parameter INVALID = 2'b00; parameter VALID = 2'b01; parameter MODIFIED = 2'b10; reg [CACHE_DATA_WID - 1 : 0] cache_var [0 : CACHE_DEPTH - 1]; reg [CACHE_TAG_randname_WID - 1 : 0] cache_randname_contr [0 : CACHE_DEPTH - 1]; reg [DATA_WID - 1 : 0] data_rand_lv5_lv5_reg; reg [DATA_WID - 1 : 0] data_rand_lv5_mem_reg; reg [31:0] zeros = 32'h0; initial begin for (i = 0; i<CACHE_DEPTH; i++) begin cache_var[i] = {CACHE_DATA_WID{1'b0}}; cache_randname_contr[i] = {CACHE_TAG_randname_WID{1'b0}}; end end assign data_rand_lv5_lv5 = data_rand_lv5_lv5_reg; assign data_rand_lv5_mem = data_rand_lv5_mem_reg; generate for(genvar gi = 1; gi<=ASSOC; gi++) begin assign cache_randname_randname[gi*randname_WID - 1 : (gi-1)*randname_WID] = cache_randname_contr[{index_randname,{ASSOC_WID{1'b0}}}+gi-1][CACHE_randname_MSB : CACHE_randname_LSB]; assign cache_randname_tag [gi*TAG_WID - 1 : (gi-1)*TAG_WID ] = cache_randname_contr[{index_randname,{ASSOC_WID{1'b0}}}+gi-1][CACHE_TAG_MSB : CACHE_TAG_LSB ]; end endgenerate always @(posedge clk) begin data_rand_lv5_lv5_reg <= 32'hz; data_rand_lv5_mem_reg <= 32'hz; addr_rand_lv5_mem <= 32'h0; data_in_rand_lv5_lv5 <= 1'bz; rand_lv5_lv5_req_lv5 <= 1'b0; mem_rd <= 1'b0; mem_wr <= 1'b0; lv5_wr_done <= 1'b0; if(lv5_rd || lv5_wr) begin if(blk_hit_randname) begin if(lv5_rd) begin if(!cp_in_cache) begin rand_lv5_lv5_req_lv5 <= 1'b1; if(rand_lv5_lv5_gnt_lv5) begin data_rand_lv5_lv5_reg <= cache_var[{index_randname,blk_access_randname}]; data_in_rand_lv5_lv5 <= 1'b1; blk_accessed_main <= blk_access_randname; end end end if(lv5_wr) begin cache_var[{index_randname,blk_access_randname}] <= data_rand_lv5_lv5; `CACHE_CURRENT_randname <= MODIFIED; blk_accessed_main <= blk_access_randname; lv5_wr_done <= 1'b1; end end else if(blk_free) begin mem_rd <= 1'b1; addr_rand_lv5_mem <= {tag_randname, index_randname, {OFFSET_WID{1'b0}}}; if(data_in_rand_lv5_mem) begin cache_var[{index_randname,blk_access_randname}] <= data_rand_lv5_mem; `CACHE_CURRENT_randname <= VALID; `CACHE_CURRENT_TAG <= tag_randname; end end else begin case(`CACHE_CURRENT_randname) VALID: `CACHE_CURRENT_randname <= INVALID; MODIFIED: begin mem_wr <= 1'b1; addr_rand_lv5_mem <= {`CACHE_CURRENT_TAG, index_randname, {OFFSET_WID{1'b0}}}; data_rand_lv5_mem_reg <= cache_var[{index_randname,blk_access_randname}]; if(mem_wr_done) begin `CACHE_CURRENT_randname <= INVALID; mem_wr <= 1'b0; addr_rand_lv5_mem <= 32'h0; data_rand_lv5_mem_reg <= 32'hz; end end default: `CACHE_CURRENT_randname <= INVALID; endcase end end end endmodule
module  flat_mod_19 #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter TAG_WID = `TAG_WID_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 , parameter INVALID = 0 )( input cmd_rd , input cmd_wr , input [TAG_MSB : TAG_LSB] tag_randname , input [ASSOC*randname_WID - 1 : 0 ] cache_randname_randname , input [ASSOC*TAG_WID - 1 : 0 ] cache_randname_tag , output reg [ASSOC - 1 : 0 ] access_blk_randname ); integer i; wire [randname_WID - 1 : 0] cache_randname [ASSOC - 1 : 0]; wire [TAG_WID - 1 : 0] cache_tag [ASSOC - 1 : 0]; generate for(genvar gi = 1; gi<=ASSOC; gi++) begin : divide assign cache_randname[gi - 1] = cache_randname_randname[gi*randname_WID - 1 : (gi-1)*randname_WID]; assign cache_tag [gi - 1] = cache_randname_tag [gi*TAG_WID - 1 : (gi-1)*TAG_WID]; end endgenerate always @* begin if(cmd_rd || cmd_wr) begin for(i = 0; i < ASSOC; i++) begin if(cache_randname[i] != INVALID && cache_tag[i] == tag_randname) access_blk_randname[i] = 1'b1; else access_blk_randname[i] = 1'b0; end end else begin for(i = 0; i < ASSOC; i++) begin access_blk_randname[i] = 1'b0; end end end endmodule
module addr_segregator_randname #( parameter ADDR_WID = `ADDR_WID_lv5 , parameter INDEX_MSB = `INDEX_MSB_lv5 , parameter INDEX_LSB = `INDEX_LSB_lv5 , parameter OFFSET_MSB = `OFFSET_MSB_lv5 , parameter OFFSET_LSB = `OFFSET_LSB_lv5 , parameter TAG_MSB = `TAG_MSB_lv5 , parameter TAG_LSB = `TAG_LSB_lv5 )( input cmd_rd , input cmd_wr , input [ADDR_WID - 1 : 0] address , output reg [INDEX_MSB : INDEX_LSB] index_randname , output reg [TAG_MSB : TAG_LSB] tag_randname , output reg [OFFSET_MSB : OFFSET_LSB] blk_offset_randname ); reg [ADDR_WID - 1 : 0] zeros = 0; always @ * begin if(cmd_rd || cmd_wr) begin index_randname = address[INDEX_MSB : INDEX_LSB]; tag_randname = address[TAG_MSB : TAG_LSB]; blk_offset_randname = address[OFFSET_MSB : OFFSET_LSB]; end else begin index_randname = zeros[INDEX_MSB : INDEX_LSB]; tag_randname = zeros[TAG_MSB : TAG_LSB]; blk_offset_randname = zeros[OFFSET_MSB : OFFSET_LSB]; end end endmodule
module  flat_mod_20 #( parameter ASSOC = `ASSOC_lv5 )( input cmd_rd , input cmd_wr , input [ASSOC - 1 : 0] access_blk_randname , output reg blk_hit_randname ); always @* begin if(cmd_rd || cmd_wr) begin if(|access_blk_randname == 1'b1) blk_hit_randname = 1'b1; else blk_hit_randname = 1'b0; end else blk_hit_randname = 1'b0; end endmodule
module blk_to_be_accessed_md #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 )( input blk_hit_randname , input [ASSOC - 1 : 0] access_blk_randname , input [ASSOC_WID - 1 : 0] lru_replacement_randname , input [ASSOC_WID - 1 : 0] free_blk_num , input blk_free , output reg [ASSOC_WID - 1 : 0] blk_access_randname ); always @* begin if(blk_hit_randname) begin blk_access_randname = 0; for(int i = 0; i < ASSOC; i++) begin if(access_blk_randname[i] == 1'b1) blk_access_randname = i; end end else if(blk_free) blk_access_randname = free_blk_num; else blk_access_randname = lru_replacement_randname; end endmodule 
module free_blk_md #( parameter ASSOC = `ASSOC_lv5 , parameter ASSOC_WID = `ASSOC_WID_lv5 , parameter randname_WID = `randname_WID_lv5 , parameter INVALID = 0 )( input blk_hit_randname , input [ASSOC*randname_WID - 1 : 0] cache_randname_randname , output reg blk_free , output reg [ASSOC_WID - 1 : 0] free_blk_num ); integer i; wire [randname_WID - 1 : 0] cache_randname [ASSOC - 1 : 0]; generate for(genvar gi = 1; gi<=ASSOC; gi++) begin : divide assign cache_randname[gi - 1] = cache_randname_randname[gi*randname_WID - 1 : (gi-1)*randname_WID]; end endgenerate always @* begin blk_free = 1'b0; free_blk_num = 0; if(blk_hit_randname == 1'b0) begin for (i = 0; i < ASSOC; i++) begin if(cache_randname[i] == INVALID) begin blk_free = 1'b1; free_blk_num = i; end end end end endmodule